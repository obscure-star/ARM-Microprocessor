-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- PROGRAM		"Quartus Prime"
-- VERSION		"Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition"
-- CREATED		"Wed Nov 24 21:02:08 2021"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Control_proc IS 
	PORT
	(
		Op :  IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		RegDst :  OUT  STD_LOGIC;
		ALUSrc :  OUT  STD_LOGIC;
		MemtoReg :  OUT  STD_LOGIC;
		RegWrite :  OUT  STD_LOGIC;
		MemRead :  OUT  STD_LOGIC;
		MemWrite :  OUT  STD_LOGIC;
		Branch :  OUT  STD_LOGIC;
		ALUOp1 :  OUT  STD_LOGIC;
		ALUOp0 :  OUT  STD_LOGIC
	);
END Control_proc;

ARCHITECTURE bdf_type OF Control_proc IS 

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;


BEGIN 
RegDst <= SYNTHESIZED_WIRE_32;
MemtoReg <= SYNTHESIZED_WIRE_31;
MemRead <= SYNTHESIZED_WIRE_31;
MemWrite <= SYNTHESIZED_WIRE_5;
Branch <= SYNTHESIZED_WIRE_29;
ALUOp1 <= SYNTHESIZED_WIRE_32;
ALUOp0 <= SYNTHESIZED_WIRE_29;



SYNTHESIZED_WIRE_30 <= SYNTHESIZED_WIRE_0 AND SYNTHESIZED_WIRE_1 AND SYNTHESIZED_WIRE_2 AND Op(3) AND SYNTHESIZED_WIRE_3 AND SYNTHESIZED_WIRE_4;


SYNTHESIZED_WIRE_1 <= NOT(Op(0));



SYNTHESIZED_WIRE_2 <= NOT(Op(1));



SYNTHESIZED_WIRE_0 <= NOT(Op(2));



SYNTHESIZED_WIRE_3 <= NOT(Op(4));



SYNTHESIZED_WIRE_4 <= NOT(Op(5));



ALUSrc <= SYNTHESIZED_WIRE_5 OR SYNTHESIZED_WIRE_30 OR SYNTHESIZED_WIRE_31;


SYNTHESIZED_WIRE_29 <= Op(2) AND SYNTHESIZED_WIRE_8 AND SYNTHESIZED_WIRE_9 AND SYNTHESIZED_WIRE_10 AND SYNTHESIZED_WIRE_11 AND SYNTHESIZED_WIRE_12;


SYNTHESIZED_WIRE_8 <= NOT(Op(0));



SYNTHESIZED_WIRE_9 <= NOT(Op(1));



SYNTHESIZED_WIRE_10 <= NOT(Op(3));



SYNTHESIZED_WIRE_11 <= NOT(Op(4));



SYNTHESIZED_WIRE_12 <= NOT(Op(5));



SYNTHESIZED_WIRE_31 <= SYNTHESIZED_WIRE_13 AND Op(0) AND Op(1) AND SYNTHESIZED_WIRE_14 AND SYNTHESIZED_WIRE_15 AND Op(5);


SYNTHESIZED_WIRE_13 <= NOT(Op(2));



SYNTHESIZED_WIRE_14 <= NOT(Op(3));



SYNTHESIZED_WIRE_15 <= NOT(Op(4));



SYNTHESIZED_WIRE_32 <= SYNTHESIZED_WIRE_16 AND SYNTHESIZED_WIRE_17 AND SYNTHESIZED_WIRE_18 AND SYNTHESIZED_WIRE_19 AND SYNTHESIZED_WIRE_20 AND SYNTHESIZED_WIRE_21;


SYNTHESIZED_WIRE_17 <= NOT(Op(0));



SYNTHESIZED_WIRE_18 <= NOT(Op(1));



SYNTHESIZED_WIRE_16 <= NOT(Op(2));



SYNTHESIZED_WIRE_19 <= NOT(Op(3));



SYNTHESIZED_WIRE_20 <= NOT(Op(4));



SYNTHESIZED_WIRE_21 <= NOT(Op(5));



RegWrite <= SYNTHESIZED_WIRE_31 OR SYNTHESIZED_WIRE_30 OR SYNTHESIZED_WIRE_32;


SYNTHESIZED_WIRE_5 <= SYNTHESIZED_WIRE_25 AND Op(0) AND Op(1) AND Op(3) AND SYNTHESIZED_WIRE_26 AND Op(5);


SYNTHESIZED_WIRE_25 <= NOT(Op(2));



SYNTHESIZED_WIRE_26 <= NOT(Op(4));



END bdf_type;